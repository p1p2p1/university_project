`timescale 1ns/1ns

module tb_calculator();

reg [5:0]   x_data;
reg [5:0]   y_data;

wire [6:0]  w_add;
wire [6:0]  w_sub;
wire [11:0] w_mul;
wire [5:0]  w_div;

initial begin
    x_data=6'd4;
    y_data=6'd2;

#10 x_data=6'd5;
    y_data=6'd6;     

#10 x_data=6'd7;
    y_data=6'd2;
end

calculator  U0_calculator(
                        .o_add  (w_add ), 
                        .o_sub  (w_sub ), 
                        .o_mul  (w_mul ), 
                        .o_div  (w_div ), 
                        .i_data1(x_data), 
                        .i_data2(y_data)
                        );
endmodule
